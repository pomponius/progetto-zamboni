LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_misc.all;

ENTITY filter IS
PORT ( CLK, RSTN, START, RD_DATA_OUT : IN STD_LOGIC;
	DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	ADDRESS_DATA_OUT : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
	DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	DONE: OUT STD_LOGIC);
END filter;

ARCHITECTURE Structural OF filter IS

COMPONENT ram
	PORT(DATA_IN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ADDRESS: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		CS, CLK, WRN, RD: IN STD_LOGIC;
		DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT register_nbit IS
	GENERIC(N: INTEGER :=8);
	PORT (R : IN STD_LOGIC_VECTOR((N-1) DOWNTO 0);
		Clk, Rstn : IN STD_LOGIC;
		Q : OUT STD_LOGIC_VECTOR((N-1) DOWNTO 0));
END COMPONENT;

COMPONENT counter_nbit IS
	GENERIC(N: INTEGER := 10);
	PORT ( Clk, Clrn, E : IN STD_LOGIC;
		COUNT : BUFFER STD_LOGIC_VECTOR((N-1) DOWNTO 0);
		MAX_VAL: OUT STD_LOGIC);
END COMPONENT;

COMPONENT subtractor_nbit IS
	GENERIC(N: INTEGER := 10);
	PORT ( A, B : IN STD_LOGIC_VECTOR((N-1) DOWNTO 0);
		DIFF: BUFFER STD_LOGIC_VECTOR((N-1) DOWNTO 0);
		OVERFLOW, UNDERFLOW, OV255, OV127, UN_256, UN_128: OUT STD_LOGIC);
END COMPONENT;

--CONTROLL SIGNALS
	--FROM CONTROL UNIT TO DATA PATH
SIGNAL RESET_ALL_N, ENABLE_COUNTER, LOAD_MEM_A_N, NEXT_VALUE, NEXT_VALUE_N, OUT_OF_RANGE, MIN_MAXN, BUSY: STD_LOGIC;
SIGNAL OPERATION: STD_LOGIC_VECTOR(1 DOWNTO 0);
	--FROM DATA PATH TO CONTROL UNIT
SIGNAL OVER255, OVER127, UNDER_256, UNDER_128, OVERFLOW, UNDERFLOW, COUNTER_OVERFLOW, SKIP: STD_LOGIC;


--BUS
SIGNAL Xn, Xn_1, Yn, Yn_1, Yn_2: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL Xn_4, Xn_1_2, Temp, Result, Yn_1_05, Yn_2_025, ADDRESS: STD_LOGIC_VECTOR(9 DOWNTO 0);

--OTHERS
SIGNAL ENABLE_CLK: STD_LOGIC;
SIGNAL OPERAND_A, OPERAND_B, ADDRESS_MEMB: STD_LOGIC_VECTOR(9 DOWNTO 0);

--CONTROL UNIT STATES
TYPE State_type IS (STANDBY, LOADING_MEMORY, OPERATION_1, OPERATION_2, OPERATION_3, ALL_DONE);
SIGNAL STATE, NEXT_STATE : State_type;

BEGIN


--DATA PATH

ENABLE_CLK<=CLK AND NEXT_VALUE;
SKIP<=nor_reduce(Yn_1_05) AND nor_reduce(Yn_2_025);

--MEMORY DECLARATION
NEXT_VALUE_N <= NOT(NEXT_VALUE);
Mem_A: ram PORT MAP(DATA_IN, ADDRESS, '1', CLK, LOAD_MEM_A_N, '1', Xn);
ADDRESS_MEMB<=ADDRESS WHEN BUSY='1' ELSE
			ADDRESS_DATA_OUT;
Mem_B: ram PORT MAP(Yn, ADDRESS_MEMB, '1', CLK, NEXT_VALUE_N, RD_DATA_OUT, DATA_OUT);

--REGISTER DECLARATION
Reg_Xn_1: register_nbit GENERIC MAP(8) PORT MAP(Xn, ENABLE_CLK, RESET_ALL_N, Xn_1);
Reg_Yn_1: register_nbit GENERIC MAP(8) PORT MAP(Yn, ENABLE_CLK, RESET_ALL_N, Yn_1);
Reg_Yn_2: register_nbit GENERIC MAP(8) PORT MAP(Yn_1, ENABLE_CLK, RESET_ALL_N, Yn_2);
Reg_Temp: register_nbit GENERIC MAP(10) PORT MAP(Result, CLK, RESET_ALL_N, Temp);

--ADDRESS COUNTER
Addr_Cont: counter_nbit GENERIC MAP(10) PORT MAP(CLK, RESET_ALL_N, ENABLE_COUNTER, ADDRESS, COUNTER_OVERFLOW);

--MOLTIPLICATION AND DIVISIONS
Xn_4<= Xn&"00";
Xn_1_2<= Xn_1(7)&Xn_1&"0";
Yn_1_05<=Yn_1(7)&Yn_1(7)&Yn_1(7)&Yn_1(7 DOWNTO 1);
Yn_2_025<=Yn_2(7)&Yn_2(7)&Yn_2(7)&Yn_2(7)&Yn_1(7 DOWNTO 2);

--ALU
OPERAND_A<=Xn_1_2 WHEN OPERATION(0)='0' ELSE
			Yn_2_025 WHEN OPERATION(1)='0' ELSE
			Yn_1_05 WHEN OPERATION (1)='1';
OPERAND_B<=Xn_4 WHEN OPERATION(0)='0' ELSE
			Temp;
Sub: subtractor_nbit GENERIC MAP(10) PORT MAP(OPERAND_A, OPERAND_B, Result, OVERFLOW, UNDERFLOW, OVER255, OVER127, UNDER_256, UNDER_128);

--RESULT
Yn<=Result(7 DOWNTO 0) WHEN OUT_OF_RANGE='0' ELSE
	"01111111" WHEN MIN_MAXN='0' ELSE
	"10000000" WHEN MIN_MAXN='1';

	
	
--CONTROL UNIT
PROCESS (STATE, START, NEXT_VALUE, COUNTER_OVERFLOW) -- state table
BEGIN
	CASE STATE IS 
		WHEN STANDBY=>
			IF(START='1') THEN
				NEXT_STATE<=LOADING_MEMORY;
			ELSE
				NEXT_STATE<=STANDBY;
			END IF;
		WHEN LOADING_MEMORY=>
			IF START='0' THEN
				NEXT_STATE<=STANDBY;
			ELSIF(COUNTER_OVERFLOW='1') THEN
				NEXT_STATE<=OPERATION_1;
			ELSE
				NEXT_STATE<=LOADING_MEMORY;
			END IF;
		WHEN OPERATION_1=>
			IF START='0' THEN
				NEXT_STATE<=STANDBY;
			ELSIF (NEXT_VALUE='1')THEN
				IF COUNTER_OVERFLOW='1' THEN
					NEXT_STATE<=ALL_DONE;
				ELSE
					NEXT_STATE<=OPERATION_1;
				END IF;
			ELSE
				NEXT_STATE<=OPERATION_2;
			END IF;
		WHEN OPERATION_2=>
			IF START='0' THEN
				NEXT_STATE<=STANDBY;
			ELSIF (NEXT_VALUE='1')THEN
				IF COUNTER_OVERFLOW='1' THEN
					NEXT_STATE<=ALL_DONE;
				ELSE
					NEXT_STATE<=OPERATION_1;
				END IF;
			ELSE
				NEXT_STATE<=OPERATION_3;
			END IF;	
		WHEN OPERATION_3=>
			IF START='0' THEN
				NEXT_STATE<=STANDBY;
			ELSIF COUNTER_OVERFLOW='1' THEN
				NEXT_STATE<=ALL_DONE;
			ELSE
				NEXT_STATE<=OPERATION_1;
			END IF;	
		WHEN ALL_DONE=>
			IF START='0' THEN
				NEXT_STATE<=STANDBY;
			ELSE
				NEXT_STATE<=ALL_DONE;
			END IF;
		WHEN OTHERS =>
			NEXT_STATE<=STANDBY;
	END CASE;
END PROCESS; -- state table


PROCESS (CLK) -- state flip-flops
BEGIN
	IF RSTN='0' THEN
		STATE<=STANDBY;
	ELSIF(CLK'EVENT AND CLK='1') THEN
		STATE<=NEXT_STATE;
	END IF;
END PROCESS;


PROCESS (STATE, OVER127, UNDER_128, OVER255, UNDER_256, OVERFLOW, UNDERFLOW, SKIP)
BEGIN
	CASE STATE IS 
		WHEN STANDBY=>
			RESET_ALL_N<='0';
			ENABLE_COUNTER<='0';
			LOAD_MEM_A_N<='1'; 
			NEXT_VALUE<='0';
			OUT_OF_RANGE<='0';
			MIN_MAXN<='0';
			BUSY<='0';
			DONE<='0';
			OPERATION<="00";
		WHEN LOADING_MEMORY=>
			RESET_ALL_N<='1';
			ENABLE_COUNTER<='1';
			LOAD_MEM_A_N<='0'; 
			NEXT_VALUE<='0';
			OUT_OF_RANGE<='0';
			MIN_MAXN<='0';
			BUSY<='1';
			DONE<='0';
			OPERATION<="00";
		WHEN OPERATION_1=>
			RESET_ALL_N<='1';
			IF (SKIP='1' OR OVERFLOW='1' OR UNDERFLOW='1' OR OVER255='1' OR UNDER_256='1') THEN
				ENABLE_COUNTER<='1';
				NEXT_VALUE<='1';
			ELSE
				ENABLE_COUNTER<='0';
				NEXT_VALUE<='0';
			END IF;
			LOAD_MEM_A_N<='1';
			IF SKIP='1' THEN				
				IF(OVER127='1' OR UNDER_128='1' OR OVERFLOW='1' OR UNDERFLOW='1') THEN
					OUT_OF_RANGE<='1';
				ELSE
					OUT_OF_RANGE<='0';
				END IF;
				IF(OVER127='1' OR OVERFLOW='1') THEN
					MIN_MAXN<='0';
				ELSIF(UNDER_128='1' OR UNDERFLOW='1') THEN
					MIN_MAXN<='1';
				END IF;
			ELSE
				IF(OVER255='1' OR UNDER_256='1' OR OVERFLOW='1' OR UNDERFLOW='1') THEN
					OUT_OF_RANGE<='1';
				ELSE
					OUT_OF_RANGE<='0';
				END IF;	
				IF(OVER255='1' OR OVERFLOW='1') THEN
					MIN_MAXN<='0';
				ELSIF(UNDER_256='1' OR UNDERFLOW='1') THEN
					MIN_MAXN<='1';
				END IF;
			END IF;
			BUSY<='1';
			DONE<='0';
			OPERATION<="00";
		WHEN OPERATION_2=>
			RESET_ALL_N<='1';
			IF (OVERFLOW='1' OR UNDERFLOW='1' OR OVER255='1' OR UNDER_256='1') THEN
				ENABLE_COUNTER<='1';
				NEXT_VALUE<='1';
			ELSE
				ENABLE_COUNTER<='0';
				NEXT_VALUE<='0';
			END IF;
			LOAD_MEM_A_N<='1';
			IF(OVERFLOW='1' OR UNDERFLOW='1' OR OVER255='1' OR UNDER_256='1') THEN
				OUT_OF_RANGE<='1';
			ELSE
				OUT_OF_RANGE<='0';
			END IF;
			IF(OVER255='1' OR OVERFLOW='1') THEN
				MIN_MAXN<='1';
			ELSIF(UNDER_256='1' OR UNDERFLOW='1') THEN
				MIN_MAXN<='0';
			END IF;
			BUSY<='1';
			DONE<='0';
			OPERATION<="01";
		WHEN OPERATION_3=>
			RESET_ALL_N<='1';
			ENABLE_COUNTER<='1';
			NEXT_VALUE<='1';
			LOAD_MEM_A_N<='1';
			IF(OVERFLOW='1' OR UNDERFLOW='1' OR OVER127='1' OR UNDER_128='1') THEN
				OUT_OF_RANGE<='1';
			ELSE
				OUT_OF_RANGE<='0';
			END IF;
			IF(OVER127='1' OR OVERFLOW='1') THEN
				MIN_MAXN<='0';
			ELSIF(UNDER_128='1' OR UNDERFLOW='1') THEN
				MIN_MAXN<='1';
			END IF;
			BUSY<='1';
			DONE<='0';
			OPERATION<="11";
		WHEN ALL_DONE=>
			RESET_ALL_N<='1';
			ENABLE_COUNTER<='0';
			NEXT_VALUE<='0';
			LOAD_MEM_A_N<='1';
			OUT_OF_RANGE<='0';	
			MIN_MAXN<='0';
			BUSY<='0';
			DONE<='1';
			OPERATION<="00";
	END CASE;

END PROCESS;



END Structural; 